--------------------------------------------------------------------------------
-- File Name: BitMapROMpkg.vhd
-- Title: BitMap ROM arrays
-- Version: 0.3
-- Date: 2016/12/19
-- Author: Miguel A. Risco Castillo
-- web page: http://sba.accesus.com
--
-- Description and Notes:
-- Package with bitmap images and character ROM for the SBA analog
-- video system.
--
--------------------------------------------------------------------------------
-- This version is released under the GNU/GLP license
-- if you use this component for your research please
-- include the appropriate credit of Author.
-- For commercial purposes request the appropriate
-- license from the author.
--------------------------------------------------------------------------------

Library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package Num16x24ROMPackage is

type TROM is Array(integer range <>,integer range <>) of std_logic_vector(7 downto 0);
type TBitRom is Array(integer range <>,integer range <>) of std_logic;

--NUMBER 16x24
constant NumDigits:integer:=16;
constant ChrW:integer:=16;
constant ChrH:integer:=24;
type TNumRom is Array(integer range <>) of std_logic_vector(0 to ChrW-1);
constant NumRom : TNumRom(0 to (NumDigits*ChrH)-1) :=(
       "0000011110000000",
       "0000111111000000",
       "0001111111100000",
       "0011100000110000",
       "0111000001111000",
       "0110000001111000",
       "1110000011111100",
       "1110000011011100",
       "1110000111011100",
       "1110000110011100",
       "1110001110011100",
       "1110001100011100",
       "1110011100011100",
       "1110011000011100",
       "1110111000011100",
       "1110110000011100",
       "1111110000011100",
       "1111100000011100",
       "0111100000011000",
       "0111000000011000",
       "0011000000110000",
       "0001111111100000",
       "0000111111000000",
       "0000011110000000",
       --
       "0000111100000000",
       "0001111100000000",
       "0011111100000000",
       "0000011100000000",
       "0000011100000000",
       "0000011100000000",
       "0000011100000000",
       "0000011100000000",
       "0000011100000000",
       "0000011100000000",
       "0000011100000000",
       "0000011100000000",
       "0000011100000000",
       "0000011100000000",
       "0000011100000000",
       "0000011100000000",
       "0000011100000000",
       "0000011100000000",
       "0000011100000000",
       "0000011100000000",
       "0000011100000000",
       "0011111111100000",
       "0011111111100000",
       "0011111111100000",
       --
       "0000111111000000",
       "0001111111100000",
       "0011111111110000",
       "0111100001111000",
       "1110000000011100",
       "1110000000011100",
       "1110000000011100",
       "0000000000011100",
       "0000000000011100",
       "0000000000111100",
       "0000000001111000",
       "0000011111110000",
       "0001111111100000",
       "0011111111000000",
       "0111100000000000",
       "1111000000000000",
       "1110000000000000",
       "1110000000000000",
       "1110000000000000",
       "1110000000000000",
       "1110000000001100",
       "1111111111111100",
       "1111111111111100",
       "0111111111110000",
       --
       "1111111111111000",
       "1111111111111100",
       "1111111111111100",
       "0000000000111100",
       "0000000000111000",
       "0000000001111000",
       "0000000011110000",
       "0000000111100000",
       "0000001111000000",
       "0000011110000000",
       "0000011110000000",
       "0000000111100000",
       "0000000011110000",
       "0000000001111000",
       "0000000000111100",
       "0000000000011100",
       "0000000000011100",
       "0000000000011100",
       "1110000000011100",
       "1110000000011100",
       "1111000000111100",
       "0111111111111000",
       "0011111111110000",
       "0001111111100000",
       --
       "0000000001100000",
       "0000000011110000",
       "0000000111110000",
       "0000000111110000",
       "0000001111110000",
       "0000001101110000",
       "0000011101110000",
       "0000011001110000",
       "0000111001110000",
       "0000110001110000",
       "0001110001110000",
       "0001100001110000",
       "0011100001110000",
       "0011000001110000",
       "0111000001110000",
       "0110000001110000",
       "1110000001110000",
       "1111111111111100",
       "1111111111111100",
       "0111111111111100",
       "0000000001110000",
       "0000000001110000",
       "0000000001110000",
       "0000000001110000",
       --
       "0111111111111000",
       "1111111111111100",
       "1111111111111100",
       "1110000000000000",
       "1110000000000000",
       "1110000000000000",
       "1110000000000000",
       "1110000000000000",
       "1110000000000000",
       "1111111111100000",
       "1111111111110000",
       "0111111111111000",
       "0000000000111100",
       "0000000000011100",
       "0000000000011100",
       "0000000000011100",
       "0000000000011100",
       "0000000000011100",
       "0000000000011100",
       "0000000000011100",
       "1110000000111000",
       "0111111111111000",
       "0011111111110000",
       "0000111111000000",
       --
       "0000000000111000",
       "0000000001111000",
       "0000000011110000",
       "0000000111100000",
       "0000001111000000",
       "0000011110000000",
       "0000111100000000",
       "0001111000000000",
       "0011110000000000",
       "0111100000000000",
       "0111111111100000",
       "1111111111110000",
       "1111111111111000",
       "1111000000111100",
       "1110000000011100",
       "1110000000011100",
       "1110000000011100",
       "1110000000011100",
       "1110000000011100",
       "1110000000011100",
       "0111000000111000",
       "0011111111111000",
       "0001111111110000",
       "0000111111000000",
       --
       "1111111111111000",
       "1111111111111100",
       "1111111111111100",
       "0000000000111100",
       "0000000000111100",
       "0000000000111000",
       "0000000001111000",
       "0000000001110000",
       "0000000011110000",
       "0000000011100000",
       "0000000111100000",
       "0000000111000000",
       "0000001111000000",
       "0000001110000000",
       "0000011110000000",
       "0000011100000000",
       "0000111100000000",
       "0000111000000000",
       "0001111000000000",
       "0001110000000000",
       "0001110000000000",
       "0001110000000000",
       "0001110000000000",
       "0001110000000000",
       --
       "0000011110000000",
       "0001111111100000",
       "0011111111110000",
       "0111000000111000",
       "1110000000011100",
       "1110000000011100",
       "1110000000011100",
       "1110000000011100",
       "1110000000011100",
       "1111000000111100",
       "0111111111111000",
       "0011111111110000",
       "0111111111111000",
       "1111000000111100",
       "1110000000011100",
       "1110000000011100",
       "1110000000011100",
       "1110000000011100",
       "1110000000011100",
       "1110000000011100",
       "0111000000111000",
       "0011111111110000",
       "0001111111100000",
       "0000011111000000",
       --
       "0000111111000000",
       "0001111111100000",
       "0011111111110000",
       "0111000000111000",
       "1110000000011100",
       "1110000000011100",
       "1110000000011100",
       "1110000000011100",
       "1110000000011100",
       "1110000000011100",
       "1111000000111100",
       "0111111111111100",
       "0011111111111100",
       "0001111111111000",
       "0000000001111000",
       "0000000011110000",
       "0000000111100000",
       "0000001111000000",
       "0000011110000000",
       "0000111100000000",
       "0001111000000000",
       "0011110000000000",
       "0111100000000000",
       "0111000000000000",
       --
       "0000001100000000",
       "0000001100000000",
       "0000011110000000",
       "0000011110000000",
       "0000111111000000",
       "0000111111000000",
       "0001111111100000",
       "0001110011100000",
       "0011110011110000",
       "0011100001110000",
       "0111100001111000",
       "0111000000111000",
       "1111000000111100",
       "1110000000011100",
       "1110000000011100",
       "1110000000011100",
       "1111111111111100",
       "1111111111111100",
       "1111111111111100",
       "1110000000011100",
       "1110000000011100",
       "1110000000011100",
       "1110000000011100",
       "1110000000011100",
       --
       "1111111111000000",
       "1111111111100000",
       "1111111111110000",
       "1110000000111000",
       "1110000000011100",
       "1110000000011100",
       "1110000000011100",
       "1110000000011100",
       "1110000000111100",
       "1110000001111000",
       "1111111111110000",
       "1111111111100000",
       "1111111111110000",
       "1110000001111000",
       "1110000000111100",
       "1110000000011100",
       "1110000000011100",
       "1110000000011100",
       "1110000000011100",
       "1110000000011100",
       "1110000000111000",
       "1111111111111000",
       "1111111111110000",
       "1111111111100000",
       --
       "0000011111000000",
       "0000111111100000",
       "0001111111110000",
       "0011110000111000",
       "0111100000011100",
       "1111000000011100",
       "1110000000011100",
       "1110000000000000",
       "1110000000000000",
       "1110000000000000",
       "1110000000000000",
       "1110000000000000",
       "1110000000000000",
       "1110000000000000",
       "1110000000000000",
       "1110000000000000",
       "1110000000000000",
       "1110000000000000",
       "1110000000011100",
       "0111000000011100",
       "0011100000111100",
       "0001111111111000",
       "0000111111110000",
       "0000011111100000",
       --
       "1111111100000000",
       "1111111110000000",
       "1111111111000000",
       "1110000111100000",
       "1110000011110000",
       "1110000001111000",
       "1110000000111100",
       "1110000000011100",
       "1110000000011100",
       "1110000000011100",
       "1110000000011100",
       "1110000000011100",
       "1110000000011100",
       "1110000000011100",
       "1110000000011100",
       "1110000000011100",
       "1110000000011100",
       "1110000000011100",
       "1110000000111100",
       "1110000001110000",
       "1110000111100000",
       "1111111111000000",
       "1111111110000000",
       "1111111100000000",
       --
       "1111111111111100",
       "1111111111111100",
       "1111111111111100",
       "1110000000000000",
       "1110000000000000",
       "1110000000000000",
       "1110000000000000",
       "1110000000000000",
       "1110000000000000",
       "1110000000000000",
       "1111111111110000",
       "1111111111110000",
       "1111111111110000",
       "1110000000000000",
       "1110000000000000",
       "1110000000000000",
       "1110000000000000",
       "1110000000000000",
       "1110000000000000",
       "1110000000000000",
       "1110000000000000",
       "1111111111111100",
       "1111111111111100",
       "1111111111111100",
       --
       "1111111111111100",
       "1111111111111100",
       "1111111111111100",
       "1110000000000000",
       "1110000000000000",
       "1110000000000000",
       "1110000000000000",
       "1110000000000000",
       "1110000000000000",
       "1110000000000000",
       "1111111111100000",
       "1111111111100000",
       "1111111111100000",
       "1110000000000000",
       "1110000000000000",
       "1110000000000000",
       "1110000000000000",
       "1110000000000000",
       "1110000000000000",
       "1110000000000000",
       "1110000000000000",
       "1110000000000000",
       "1110000000000000",
       "1110000000000000"
);

  function NumPx(X,Y:integer;N:unsigned) return std_logic;


end Num16x24ROMPackage;

package body Num16x24ROMPackage is

  function NumPx(X,Y:integer;N:unsigned) return std_logic is
  variable posX:integer range 0 to N'length/4-1;
  variable tmp:integer range 0 to 15;
  variable trow:std_logic_vector(0 to ChrW-1);
  begin
    posX:= N'length/4 - (X/ChrW) - 1;
    tmp := to_integer(N(4*posX+3 downto 4*posX));
    trow:= NumRom((tmp * ChrH)+Y);
    return trow(X mod ChrW);
  end;

end Num16x24ROMPackage;
