--------------------------------------------------------------------------------
-- File Name: Txt16x19ROMpkg.vhd
-- Title: Text BitMap ROM
-- Version: 0.2
-- Date: 2016/12/19
-- Author: Miguel A. Risco Castillo
-- web page: http://sba.accesus.com
--
-- Description and Notes:
-- Package with bitmap character ROM for the SBA analog
-- video system.
--
--------------------------------------------------------------------------------
-- This version is released under the GNU/GLP license
-- if you use this component for your research please
-- include the appropriate credit of Author.
-- For commercial purposes request the appropriate
-- license from the author.
--------------------------------------------------------------------------------

Library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package Txt16x19ROMPackage is

--entity TxtROM is
--    Generic (TextRom:TBitRom:=Text16x19Rom);
--    Port ( -- SBA interface
--           CLK_I : in STD_LOGIC;
--           --TxtROM interface
--           addr  : in integer range TextRom'range;
--           data  : out std_logic_vector;
--         );
--end TxtROM;


--NUMBER 16x19 "ABCDEFGHIJKLMNOPQRSTUVWXYZ #,-./:=|°"
constant NumChars:integer:=36;
constant ChrW:integer:=16;
constant ChrH:integer:=19;
type TTextRom is Array(integer range <>) of std_logic_vector(0 to ChrW-1);
constant TextRom : TTextRom(0 to (NumChars*ChrH)-1) :=(
       "0000001110000000",
       "0000011111000000",
       "0000011011000000",
       "0000011011000000",
       "0000111011100000",
       "0000110001100000",
       "0000110001100000",
       "0001110001110000",
       "0001100000110000",
       "0001100000110000",
       "0011100000111000",
       "0011000000111000",
       "0011000000011000",
       "0111111111111100",
       "0111111111111100",
       "0110000000001100",
       "1110000000001110",
       "1110000000001110",
       "1100000000000110",
       --
       "0011111111000000",
       "0011111111110000",
       "0011100001111000",
       "0011100000111000",
       "0011100000111000",
       "0011100000111000",
       "0011100000111000",
       "0011100001110000",
       "0011111111100000",
       "0011111111110000",
       "0011100001111000",
       "0011100000011100",
       "0011100000011100",
       "0011100000011100",
       "0011100000011100",
       "0011100000011100",
       "0011100000111000",
       "0011111111110000",
       "0011111111000000",
       --
       "0000001111111000",
       "0000111111111100",
       "0001111000000100",
       "0001110000000000",
       "0011100000000000",
       "0011100000000000",
       "0111000000000000",
       "0111000000000000",
       "0111000000000000",
       "0111000000000000",
       "0111000000000000",
       "0111000000000000",
       "0111000000000000",
       "0111100000000000",
       "0011100000000000",
       "0011110000000000",
       "0001111000000100",
       "0000111111111100",
       "0000001111111000",
       --
       "0011111111100000",
       "0011111111111000",
       "0011100000111100",
       "0011100000011110",
       "0011100000001110",
       "0011100000000111",
       "0011100000000111",
       "0011100000000111",
       "0011100000000111",
       "0011100000000111",
       "0011100000000111",
       "0011100000000111",
       "0011100000000111",
       "0011100000001110",
       "0011100000001110",
       "0011100000011100",
       "0011100000111100",
       "0011111111110000",
       "0011111111000000",
       --
       "0001111111111100",
       "0001111111111100",
       "0001110000000000",
       "0001110000000000",
       "0001110000000000",
       "0001110000000000",
       "0001110000000000",
       "0001110000000000",
       "0001111111111100",
       "0001111111111100",
       "0001110000000000",
       "0001110000000000",
       "0001110000000000",
       "0001110000000000",
       "0001110000000000",
       "0001110000000000",
       "0001110000000000",
       "0001111111111100",
       "0001111111111100",
       --
       "0001111111111000",
       "0001111111111000",
       "0001110000000000",
       "0001110000000000",
       "0001110000000000",
       "0001110000000000",
       "0001110000000000",
       "0001110000000000",
       "0001110000000000",
       "0001111111111000",
       "0001111111111000",
       "0001110000000000",
       "0001110000000000",
       "0001110000000000",
       "0001110000000000",
       "0001110000000000",
       "0001110000000000",
       "0001110000000000",
       "0001110000000000",
       --
       "0000000111111100",
       "0000011111111110",
       "0000111100000010",
       "0001110000000000",
       "0011100000000000",
       "0011100000000000",
       "0111000000000000",
       "0111000000000000",
       "0111000000000000",
       "0111000011111110",
       "0111000011111110",
       "0111000000001110",
       "0111000000001110",
       "0011100000001110",
       "0011100000001110",
       "0011110000001110",
       "0001111000001110",
       "0000111111111110",
       "0000001111111000",
       --
       "0011100000011100",
       "0011100000011100",
       "0011100000011100",
       "0011100000011100",
       "0011100000011100",
       "0011100000011100",
       "0011100000011100",
       "0011100000011100",
       "0011111111111100",
       "0011111111111100",
       "0011100000011100",
       "0011100000011100",
       "0011100000011100",
       "0011100000011100",
       "0011100000011100",
       "0011100000011100",
       "0011100000011100",
       "0011100000011100",
       "0011100000011100",
       --
       "0001111111111100",
       "0001111111111100",
       "0000000111000000",
       "0000000111000000",
       "0000000111000000",
       "0000000111000000",
       "0000000111000000",
       "0000000111000000",
       "0000000111000000",
       "0000000111000000",
       "0000000111000000",
       "0000000111000000",
       "0000000111000000",
       "0000000111000000",
       "0000000111000000",
       "0000000111000000",
       "0000000111000000",
       "0001111111111100",
       "0001111111111100",
       --
       "0001111111111000",
       "0001111111111000",
       "0000000000111000",
       "0000000000111000",
       "0000000000111000",
       "0000000000111000",
       "0000000000111000",
       "0000000000111000",
       "0000000000111000",
       "0000000000111000",
       "0000000000111000",
       "0000000000111000",
       "0000000000111000",
       "0000000000111000",
       "0000000000111000",
       "0000000000111000",
       "0001000001110000",
       "0001111111100000",
       "0000111111000000",
       --
       "0011100000001110",
       "0011100000011100",
       "0011100000111000",
       "0011100001110000",
       "0011100001100000",
       "0011100011100000",
       "0011100111000000",
       "0011101110000000",
       "0011101100000000",
       "0011111100000000",
       "0011101100000000",
       "0011101110000000",
       "0011100111000000",
       "0011100011100000",
       "0011100001110000",
       "0011100001110000",
       "0011100000111000",
       "0011100000011100",
       "0011100000001110",
       --
       "0001110000000000",
       "0001110000000000",
       "0001110000000000",
       "0001110000000000",
       "0001110000000000",
       "0001110000000000",
       "0001110000000000",
       "0001110000000000",
       "0001110000000000",
       "0001110000000000",
       "0001110000000000",
       "0001110000000000",
       "0001110000000000",
       "0001110000000000",
       "0001110000000000",
       "0001110000000000",
       "0001110000000000",
       "0001111111111100",
       "0001111111111100",
       --
       "0111100000011110",
       "0111100000011110",
       "0111100000011110",
       "0110110000110110",
       "0110110000110110",
       "0110110000100110",
       "0110011001100110",
       "0110011001100110",
       "0110011001000110",
       "0110001111000110",
       "0110001111000110",
       "0110000110000110",
       "0110000110000110",
       "0110000000000110",
       "0110000000000110",
       "0110000000000110",
       "0110000000000110",
       "0110000000000110",
       "0110000000000110",
       --
       "0011110000011100",
       "0011110000011100",
       "0011111000011100",
       "0011111000011100",
       "0011111000011100",
       "0011101100011100",
       "0011101100011100",
       "0011101100011100",
       "0011100110011100",
       "0011100110011100",
       "0011100110011100",
       "0011100011011100",
       "0011100011011100",
       "0011100011011100",
       "0011100001111100",
       "0011100001111100",
       "0011100001111100",
       "0011100000111100",
       "0011100000111100",
       --
       "0000001111100000",
       "0000111111110000",
       "0001110000111000",
       "0011100000011100",
       "0011100000011100",
       "0011000000001110",
       "0111000000001110",
       "0111000000001110",
       "0111000000001110",
       "0111000000001110",
       "0111000000001110",
       "0111000000001110",
       "0111000000001110",
       "0111000000001100",
       "0011100000011100",
       "0011100000011100",
       "0001110000111000",
       "0000111111110000",
       "0000011111000000",
       --
       "0011111111100000",
       "0011111111111000",
       "0011100000111100",
       "0011100000011110",
       "0011100000001110",
       "0011100000001110",
       "0011100000001110",
       "0011100000001110",
       "0011100000011100",
       "0011100000111100",
       "0011111111111000",
       "0011111111100000",
       "0011100000000000",
       "0011100000000000",
       "0011100000000000",
       "0011100000000000",
       "0011100000000000",
       "0011100000000000",
       "0011100000000000",
       --
       "0000001111110000",
       "0000111111111000",
       "0001111000111100",
       "0011110000001110",
       "0011100000001110",
       "0011100000000111",
       "0111000000000111",
       "0111000000000111",
       "0111000000000111",
       "0111000000000111",
       "0111000000000111",
       "0111000000000111",
       "0111000011000111",
       "0111000011100110",
       "0011100001110110",
       "0011100000111110",
       "0001111000011100",
       "0000111111111110",
       "0000011111100110",
       --
       "0011111111000000",
       "0011111111110000",
       "0011100001111000",
       "0011100000111000",
       "0011100000111000",
       "0011100000111000",
       "0011100000111000",
       "0011100001110000",
       "0011111111100000",
       "0011111110000000",
       "0011100011000000",
       "0011100011100000",
       "0011100001100000",
       "0011100001110000",
       "0011100000110000",
       "0011100000111000",
       "0011100000111000",
       "0011100000011000",
       "0011100000011100",
       --
       "0000001111111000",
       "0000111111111100",
       "0001111000000100",
       "0011100000000000",
       "0011100000000000",
       "0011100000000000",
       "0011110000000000",
       "0001111000000000",
       "0000111111000000",
       "0000011111110000",
       "0000000011111100",
       "0000000000111100",
       "0000000000011110",
       "0000000000001110",
       "0000000000001110",
       "0000000000001110",
       "0010000000111100",
       "0011111111111000",
       "0000111111100000",
       --
       "0011111111111110",
       "0011111111111110",
       "0000000111000000",
       "0000000111000000",
       "0000000111000000",
       "0000000111000000",
       "0000000111000000",
       "0000000111000000",
       "0000000111000000",
       "0000000111000000",
       "0000000111000000",
       "0000000111000000",
       "0000000111000000",
       "0000000111000000",
       "0000000111000000",
       "0000000111000000",
       "0000000111000000",
       "0000000111000000",
       "0000000111000000",
       --
       "0011100000001110",
       "0011100000001110",
       "0011100000001110",
       "0011100000001110",
       "0011100000001110",
       "0011100000001110",
       "0011100000001110",
       "0011100000001110",
       "0011100000001110",
       "0011100000001110",
       "0011100000001110",
       "0011100000001110",
       "0011100000001110",
       "0011100000001110",
       "0011100000001110",
       "0011110000011100",
       "0001110000111100",
       "0000111111111000",
       "0000011111100000",
       --
       "0111000000000011",
       "0111000000000111",
       "0111000000000111",
       "0011000000000110",
       "0011100000001110",
       "0011100000001110",
       "0001100000001100",
       "0001110000011100",
       "0001110000011100",
       "0000110000011000",
       "0000111000111000",
       "0000111000111000",
       "0000011000110000",
       "0000011101110000",
       "0000011101110000",
       "0000001101100000",
       "0000001101100000",
       "0000001111100000",
       "0000000111000000",
       --
       "0111000000001110",
       "0111000000001110",
       "0111000000001110",
       "0111000000001110",
       "0111000000001110",
       "0111000000001110",
       "0111000110001110",
       "0111000110001110",
       "0111001111001110",
       "0111001111001110",
       "0011001111001100",
       "0011001001101100",
       "0011011001101100",
       "0011011001101100",
       "0011010000111100",
       "0011110000111100",
       "0011110000111100",
       "0011100000011100",
       "0011100000011100",
       --
       "0111000000001110",
       "0011100000011100",
       "0001100000011000",
       "0001110000111000",
       "0000111001110000",
       "0000111001110000",
       "0000011111100000",
       "0000001111000000",
       "0000001111000000",
       "0000001111000000",
       "0000011111000000",
       "0000011111100000",
       "0000111001110000",
       "0000111001110000",
       "0001110000111000",
       "0011100000011100",
       "0011100000011100",
       "0111000000001110",
       "1110000000000111",
       --
       "1110000000000011",
       "0111000000000111",
       "0111100000000111",
       "0011100000001110",
       "0001110000011100",
       "0001110000011100",
       "0000111000111000",
       "0000111000111000",
       "0000011101110000",
       "0000001111100000",
       "0000001111100000",
       "0000000111000000",
       "0000000111000000",
       "0000000111000000",
       "0000000111000000",
       "0000000111000000",
       "0000000111000000",
       "0000000111000000",
       "0000000111000000",
       --
       "1011111111111100",
       "0011111111111100",
       "0000000000001100",
       "0000000000011100",
       "0000000000111000",
       "0000000000110000",
       "0000000001110000",
       "0000000011100000",
       "0000000011000000",
       "0000000111000000",
       "0000000110000000",
       "0000001110000000",
       "0000011100000000",
       "0000011000000000",
       "0000111000000000",
       "0000110000000000",
       "0001100000000000",
       "0011111111111100",
       "0011111111111100",
       --
       "0000000000000000",
       "0000000000000000",
       "0000000000000000",
       "0000000000000000",
       "0000000000000000",
       "0000000000000000",
       "0000000000000000",
       "0000000000000000",
       "0000000000000000",
       "0000000000000000",
       "0000000000000000",
       "0000000000000000",
       "0000000000000000",
       "0000000000000000",
       "0000000000000000",
       "0000000000000000",
       "0000000000000000",
       "0000000000000000",
       "0000000000000000",
       --
       "0000000110011000",
       "0000000110011000",
       "0000000110011000",
       "0000001100110000",
       "0000001100110000",
       "0011111111111111",
       "0011111111111111",
       "0000001100110000",
       "0000001100110000",
       "0000001100110000",
       "0000011001100000",
       "0000011001100000",
       "0111111111111110",
       "0111111111111110",
       "0000011001100000",
       "0000011001100000",
       "0000111011100000",
       "0000110011000000",
       "0000110011000000",
       --
       "0000000000000000",
       "0000000000000000",
       "0000000000000000",
       "0000000000000000",
       "0000000000000000",
       "0000000000000000",
       "0000000000000000",
       "0000000000000000",
       "0000000000000000",
       "0000000000000000",
       "0000000111000000",
       "0000001111100000",
       "0000001111100000",
       "0000000111100000",
       "0000000111100000",
       "0000000111100000",
       "0000001111000000",
       "0000011110000000",
       "0000111000000000",
       --
       "0000000000000000",
       "0000000000000000",
       "0000000000000000",
       "0000000000000000",
       "0000000000000000",
       "0000000000000000",
       "0000000000000000",
       "0000000000000000",
       "0000000000000000",
       "0000111111110000",
       "0000111111110000",
       "0000000000000000",
       "0000000000000000",
       "0000000000000000",
       "0000000000000000",
       "0000000000000000",
       "0000000000000000",
       "0000000000000000",
       "0000000000000000",
       --
       "0000000000000000",
       "0000000000000000",
       "0000000000000000",
       "0000000000000000",
       "0000000000000000",
       "0000000000000000",
       "0000000000000000",
       "0000000000000000",
       "0000000000000000",
       "0000000000000000",
       "0000000000000000",
       "0000000000000000",
       "0000000000000000",
       "0000000000000000",
       "0000000111000000",
       "0000001111100000",
       "0000001111100000",
       "0000001111100000",
       "0000000111000000",
       --
       "0000000000011100",
       "0000000000011000",
       "0000000000111000",
       "0000000000110000",
       "0000000000110000",
       "0000000001110000",
       "0000000001100000",
       "0000000011100000",
       "0000000011000000",
       "0000000111000000",
       "0000000110000000",
       "0000000110000000",
       "0000001100000000",
       "0000001100000000",
       "0000011100000000",
       "0000011000000000",
       "0000111000000000",
       "0000110000000000",
       "0000110000000000",
       --
       "0000000000000000",
       "0000000000000000",
       "0000000000000000",
       "0000000110000000",
       "0000001111000000",
       "0000001111000000",
       "0000000110000000",
       "0000000000000000",
       "0000000000000000",
       "0000000000000000",
       "0000000000000000",
       "0000000000000000",
       "0000000000000000",
       "0000000110000000",
       "0000001111000000",
       "0000001111000000",
       "0000000110000000",
       "0000000000000000",
       "0000000000000000",
       --
       "0000000000000000",
       "0000000000000000",
       "0000000000000000",
       "0000000000000000",
       "0000000000000000",
       "0000000000000000",
       "0011111111111100",
       "0011111111111100",
       "0000000000000000",
       "0000000000000000",
       "0000000000000000",
       "0011111111111100",
       "0011111111111100",
       "0000000000000000",
       "0000000000000000",
       "0000000000000000",
       "0000000000000000",
       "0000000000000000",
       "0000000000000000",
       --
       "0000000111000000",
       "0000000111000000",
       "0000000111000000",
       "0000000111000000",
       "0000000111000000",
       "0000000111000000",
       "0000000111000000",
       "0000000111000000",
       "0000000111000000",
       "0000000111000000",
       "0000000111000000",
       "0000000111000000",
       "0000000111000000",
       "0000000111000000",
       "0000000111000000",
       "0000000111000000",
       "0000000111000000",
       "0000000111000000",
       "0000000111000000",
       --
       "0000011111000000",
       "0000111111110000",
       "0001110001110000",
       "0011100000111000",
       "0011100000111000",
       "0011100000111000",
       "0011100000111000",
       "0001110001110000",
       "0001111111100000",
       "0000011111000000",
       "0000000000000000",
       "0000000000000000",
       "0000000000000000",
       "0000000000000000",
       "0000000000000000",
       "0000000000000000",
       "0000000000000000",
       "0000000000000000",
       "0000000000000000"
       );

  function StrPx(X,Y:integer;TextString:String) return std_logic;

end Txt16x19ROMPackage;

package body Txt16x19ROMPackage is

  function StrPx(X,Y:integer;TextString:String) return std_logic is
  variable posX:integer range 1 to TextString'length;
  variable tmp:integer range 0 to 255;
  variable trow:std_logic_vector(0 to ChrW-1);
  begin
    posX := (X/ChrW)+1;
    case character'pos(TextString(PosX)) is
      when 32 => tmp:=26;  -- ' '
      when 35 => tmp:=27;  -- '#'
      when 44 => tmp:=28;  -- ','
      when 45 => tmp:=29;  -- '-'
      when 46 => tmp:=30;  -- '.'
      when 47 => tmp:=31;  -- '/'
      when 58 => tmp:=32;  -- ':'
      when 61 => tmp:=33;  -- '='
      when 124 => tmp:=34; -- '|'
      when 176 => tmp:=35; -- '°'
      when 65 to 90  => tmp:=character'pos(TextString(PosX))-65;  -- A..Z
      when 97 to 122 => tmp:=character'pos(TextString(PosX))-97;  -- a..z
      when others => tmp := 0;
    end case;
    trow:=TextRom((tmp * ChrH)+Y);
    return trow(X mod ChrW);
  end;

end Txt16x19ROMPackage;
